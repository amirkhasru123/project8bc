module forEx;
	integer i=0;
	initial begin
		for(i=0;i<2;i++) begin
			$display("I like coding a lot");
		end
	end
endmodule
