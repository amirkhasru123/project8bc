module foreverEx;
	initial begin
		forever begin
			$display("I am done");
		end
	end
endmodule
