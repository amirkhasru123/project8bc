module random;
	initial begin
		if($random)
			$display("amir is tired and bored.");
	end
endmodule
