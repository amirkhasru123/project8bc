module forEx;
	integer i=0;
	initial begin
		for(i=0;i<10;i++)
			$display("I like coding a lot");
	end
endmodule
