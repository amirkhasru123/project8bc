module foreverEx;
	initial begin
		forever
			$display("I am done");
	end
endmodule
