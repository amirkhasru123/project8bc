module repeatEx;
	initial begin
		repeat(3) begin
			$display("I love coding");
		end
	end
endmodule
