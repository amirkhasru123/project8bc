module comment;
	initial begin
		$display("Boom"); //This comment will not be outputed
		$finish;

		/*We are doing well
		* & very excited about Verilog.
		* Thank you, Rabiul Sir for instructions.
		* */
	end
endmodule
