`define amir 1

module defineEx;
    initial begin
        if (`amir) begin
            $display("I am amir");
        end
    end
endmodule

