//In verilog double slash indicates comments. Comments are left off during the execution of code.
//
//We are dealing with come circuit blocks. So we need a module. The name of the module is counter.
module counter;
	//The module doesn't have any port_lists.
endmodule
//If we run this code, we'll get nothing as output.
