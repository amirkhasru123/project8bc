`include "define.v"

module includeEx;
	initial begin
	end
endmodule
